
module PC(
	input logic clk,
	input logic rst,
	input logic [31:0] pc_next,
	output logic [31:0] pc
);

always_ff @(posedge clk or posedge rst) begin
	if(rst)begin
		pc <= 32'h0000_0000;
	end
	else begin
		pc <= pc_next;
	end
end

endmodule