// hello there , how are you 